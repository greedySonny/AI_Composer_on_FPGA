


`define CMD_NONE                    0
`define CMD_LOAD_EMBEDDING          1
`define CMD_LOAD_ZEMBEDDING         2
`define CMD_LOAD_BIAS               3
`define CMD_LOAD_WEIGHT_I           4
`define CMD_LOAD_WEIGHT_H           5
`define CMD_LOAD_RESULT             6

`define CMD_LOAD_SIGMOID		    8
`define CMD_LOAD_TANH			    9
`define CMD_STORE_R                 10
`define CMD_STORE_Z                 11
`define CMD_LOAD_R				    12
`define CMD_STORE_H 			    13
`define CMD_STORE_LAYER 		    14
`define CMD_LOAD_LAYER			    15
`define CMD_LOAD_Z				    16
`define CMD_LOAD_H				    17
`define CMD_LOAD_ZMINUS			    18
`define CMD_INIT_H				    19
`define CMD_EXP					    20
`define CMD_ADD                     22



`define CMD_DEBUG                     25
`define CMD_LOAD_TEST			      26


